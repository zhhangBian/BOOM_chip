`include "a_defines.svh"

module mdu_diver (
  input   wire    clk,
  input   wire    rst_n,
  input   wire    flush,

  

  handshake_if.receiver receiver,
  handshake_if.sender   sender
);




endmodule