`ifndef _BOOM_PARAM_HEAD
`define _BOOM_PARAM_HEAD

`endif