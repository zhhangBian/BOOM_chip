
module e_alu(
  input   logic [31:0] r0_i;
);
  
endmodule