`inclulde "define.svh"