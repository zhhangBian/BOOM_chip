`include "a_defines.svh"

module icache #(
     
) (

)

endmodule