`include "a_defines.svh"

module storebuffer #(

) (

)



endmodule