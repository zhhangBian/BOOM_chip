

module cdb #() (
    input clk,
    input rst_n,
    input flush
);
    
endmodule