`ifndef _BOOM_CSR_HEAD
`define _BOOM_CSR_HEAD

`endif