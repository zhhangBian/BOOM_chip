`ifndef _BOOM_EXCEPTION_HEAD
`deifne _BOOM_EXCEPTION_HEAD

`define 


`endif