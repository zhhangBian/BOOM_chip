`ifndef _BOOM_DECODER_HEAD
`define _BOOM_DECODER_HEAD

`endif