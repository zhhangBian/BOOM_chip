`include "a_defines.svh"

module test #(
    parameter type T = logic[31:0]
)  (
    input logic clk,
    input logic rst_n
);




endmodule