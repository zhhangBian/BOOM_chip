`ifndef _a_iq_defines
`define _a_iq_defines

`endif