`ifndef _BOOM_EXCEPTION_HEAD
`define _BOOM_EXCEPTION_HEAD

`define 


`endif