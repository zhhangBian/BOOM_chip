`include "a_defines.svh"

module dcache #(

) (
    
)

endmodule