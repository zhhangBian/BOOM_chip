`ifndef _BOOM_HEAD
`define _BOOM_HEAD

//`define _VERILATOR
// `define _ASIC
`define _FPGA

`deifne _DIFFTEST


`include "a_macros.svh"
`include "a_csr.svh"
`include "a_mmu_defines.svh"
`include "a_structure.svh"
`include "a_interface.svh"
`include "a_alu_defines.svh"
`include "a_mdu_defines.svh"
`include "a_exception_defines.svh"

`endif
