`include "a_defines.svh"

module mmu #(

) (

)

endmodule