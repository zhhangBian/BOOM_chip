`ifndef _BOOM_HEAD
`define _BOOM_HEAD

// `define _VERILATOR
// `define _ASIC
// `define _FPGA


`include "a_params.svh"
`include "a_decoder.svh"
// `include "a_macros.svh"
`include "a_structure.svh"
`include "a_csr.svh"
`include "a_interface.svh"

`endif
