`ifndef _BOOM_MACROS_HEAD
`define _BOOM_MACROS_HEAD

`define ARF_WIDTH 5
`define ROB_WIDTH 6

`define ALU_TYPE   'd1
`define MDU_TYPE   'd2
`define LSU_TYPE   'd3
`define RESERVE    'd0

`endif
